
module img_ram (
	input clk,
	input reset,
	input [127:0] dw,
	input [7:0] addr_w,
	input write,
	input read,
	input [9:0] addr_r,
	output [7:0] dr
);

logic [7:0] m [1023:0];

assign dr = read ? m[addr_r] : 0;

//m
always_ff @(posedge clk) begin
	if(!reset) begin
		if(write) begin
			m[addr_w*16] <= dw[7:0];
			m[addr_w*16+1] <= dw[15:8];
			m[addr_w*16+2] <= dw[23:16];
			m[addr_w*16+3] <= dw[31:24];
			m[addr_w*16+4] <= dw[39:32];
			m[addr_w*16+5] <= dw[47:40];
			m[addr_w*16+6] <= dw[55:48];
			m[addr_w*16+7] <= dw[63:56];
			m[addr_w*16+8] <= dw[71:64];
			m[addr_w*16+9] <= dw[79:72];
			m[addr_w*16+10] <= dw[87:80];
			m[addr_w*16+11] <= dw[95:88];
			m[addr_w*16+12] <= dw[103:96];
			m[addr_w*16+13] <= dw[111:104];
			m[addr_w*16+14] <= dw[119:112];
			m[addr_w*16+15] <= dw[127:120];
		end
	end else begin
m[0] <= 0;
m[1] <= 0;
m[2] <= 0;
m[3] <= 0;
m[4] <= 0;
m[5] <= 0;
m[6] <= 0;
m[7] <= 0;
m[8] <= 0;
m[9] <= 0;
m[10] <= 0;
m[11] <= 0;
m[12] <= 0;
m[13] <= 0;
m[14] <= 0;
m[15] <= 0;
m[16] <= 0;
m[17] <= 0;
m[18] <= 0;
m[19] <= 0;
m[20] <= 0;
m[21] <= 0;
m[22] <= 0;
m[23] <= 0;
m[24] <= 0;
m[25] <= 0;
m[26] <= 0;
m[27] <= 0;
m[28] <= 0;
m[29] <= 0;
m[30] <= 0;
m[31] <= 0;
m[32] <= 0;
m[33] <= 0;
m[34] <= 0;
m[35] <= 0;
m[36] <= 0;
m[37] <= 0;
m[38] <= 0;
m[39] <= 0;
m[40] <= 0;
m[41] <= 0;
m[42] <= 0;
m[43] <= 0;
m[44] <= 0;
m[45] <= 0;
m[46] <= 0;
m[47] <= 0;
m[48] <= 0;
m[49] <= 0;
m[50] <= 0;
m[51] <= 0;
m[52] <= 0;
m[53] <= 0;
m[54] <= 0;
m[55] <= 0;
m[56] <= 0;
m[57] <= 0;
m[58] <= 0;
m[59] <= 0;
m[60] <= 0;
m[61] <= 0;
m[62] <= 0;
m[63] <= 0;
m[64] <= 0;
m[65] <= 0;
m[66] <= 0;
m[67] <= 0;
m[68] <= 0;
m[69] <= 0;
m[70] <= 0;
m[71] <= 0;
m[72] <= 0;
m[73] <= 0;
m[74] <= 0;
m[75] <= 0;
m[76] <= 0;
m[77] <= 0;
m[78] <= 0;
m[79] <= 0;
m[80] <= 0;
m[81] <= 0;
m[82] <= 0;
m[83] <= 0;
m[84] <= 0;
m[85] <= 0;
m[86] <= 0;
m[87] <= 0;
m[88] <= 0;
m[89] <= 0;
m[90] <= 0;
m[91] <= 0;
m[92] <= 0;
m[93] <= 0;
m[94] <= 0;
m[95] <= 0;
m[96] <= 0;
m[97] <= 0;
m[98] <= 0;
m[99] <= 0;
m[100] <= 0;
m[101] <= 0;
m[102] <= 0;
m[103] <= 0;
m[104] <= 0;
m[105] <= 0;
m[106] <= 0;
m[107] <= 0;
m[108] <= 0;
m[109] <= 0;
m[110] <= 0;
m[111] <= 0;
m[112] <= 0;
m[113] <= 0;
m[114] <= 0;
m[115] <= 0;
m[116] <= 0;
m[117] <= 0;
m[118] <= 0;
m[119] <= 0;
m[120] <= 0;
m[121] <= 0;
m[122] <= 0;
m[123] <= 0;
m[124] <= 0;
m[125] <= 0;
m[126] <= 0;
m[127] <= 0;
m[128] <= 0;
m[129] <= 0;
m[130] <= 0;
m[131] <= 0;
m[132] <= 0;
m[133] <= 0;
m[134] <= 0;
m[135] <= 0;
m[136] <= 0;
m[137] <= 0;
m[138] <= 0;
m[139] <= 0;
m[140] <= 0;
m[141] <= 0;
m[142] <= 0;
m[143] <= 0;
m[144] <= 0;
m[145] <= 0;
m[146] <= 0;
m[147] <= 0;
m[148] <= 0;
m[149] <= 0;
m[150] <= 0;
m[151] <= 0;
m[152] <= 0;
m[153] <= 0;
m[154] <= 0;
m[155] <= 0;
m[156] <= 0;
m[157] <= 0;
m[158] <= 0;
m[159] <= 0;
m[160] <= 0;
m[161] <= 0;
m[162] <= 0;
m[163] <= 0;
m[164] <= 0;
m[165] <= 0;
m[166] <= 0;
m[167] <= 0;
m[168] <= 0;
m[169] <= 0;
m[170] <= 0;
m[171] <= 0;
m[172] <= 0;
m[173] <= 0;
m[174] <= 0;
m[175] <= 0;
m[176] <= 0;
m[177] <= 0;
m[178] <= 0;
m[179] <= 0;
m[180] <= 0;
m[181] <= 0;
m[182] <= 0;
m[183] <= 0;
m[184] <= 0;
m[185] <= 0;
m[186] <= 0;
m[187] <= 0;
m[188] <= 0;
m[189] <= 0;
m[190] <= 0;
m[191] <= 0;
m[192] <= 0;
m[193] <= 0;
m[194] <= 0;
m[195] <= 0;
m[196] <= 0;
m[197] <= 0;
m[198] <= 0;
m[199] <= 0;
m[200] <= 0;
m[201] <= 0;
m[202] <= 0;
m[203] <= 0;
m[204] <= 0;
m[205] <= 0;
m[206] <= 0;
m[207] <= 0;
m[208] <= 0;
m[209] <= 0;
m[210] <= 0;
m[211] <= 0;
m[212] <= 0;
m[213] <= 0;
m[214] <= 0;
m[215] <= 0;
m[216] <= 0;
m[217] <= 0;
m[218] <= 0;
m[219] <= 0;
m[220] <= 0;
m[221] <= 0;
m[222] <= 0;
m[223] <= 0;
m[224] <= 0;
m[225] <= 0;
m[226] <= 0;
m[227] <= 0;
m[228] <= 0;
m[229] <= 0;
m[230] <= 0;
m[231] <= 0;
m[232] <= 0;
m[233] <= 0;
m[234] <= 0;
m[235] <= 0;
m[236] <= 0;
m[237] <= 0;
m[238] <= 0;
m[239] <= 0;
m[240] <= 0;
m[241] <= 0;
m[242] <= 0;
m[243] <= 0;
m[244] <= 0;
m[245] <= 0;
m[246] <= 0;
m[247] <= 0;
m[248] <= 0;
m[249] <= 0;
m[250] <= 0;
m[251] <= 0;
m[252] <= 0;
m[253] <= 0;
m[254] <= 0;
m[255] <= 0;
m[256] <= 0;
m[257] <= 0;
m[258] <= 0;
m[259] <= 0;
m[260] <= 0;
m[261] <= 0;
m[262] <= 0;
m[263] <= 0;
m[264] <= 0;
m[265] <= 0;
m[266] <= 0;
m[267] <= 0;
m[268] <= 0;
m[269] <= 0;
m[270] <= 0;
m[271] <= 0;
m[272] <= 0;
m[273] <= 0;
m[274] <= 0;
m[275] <= 0;
m[276] <= 0;
m[277] <= 0;
m[278] <= 0;
m[279] <= 0;
m[280] <= 0;
m[281] <= 0;
m[282] <= 0;
m[283] <= 0;
m[284] <= 0;
m[285] <= 0;
m[286] <= 0;
m[287] <= 0;
m[288] <= 0;
m[289] <= 0;
m[290] <= 0;
m[291] <= 0;
m[292] <= 0;
m[293] <= 0;
m[294] <= 0;
m[295] <= 0;
m[296] <= 0;
m[297] <= 0;
m[298] <= 0;
m[299] <= 0;
m[300] <= 0;
m[301] <= 0;
m[302] <= 0;
m[303] <= 0;
m[304] <= 0;
m[305] <= 0;
m[306] <= 0;
m[307] <= 0;
m[308] <= 0;
m[309] <= 0;
m[310] <= 0;
m[311] <= 0;
m[312] <= 0;
m[313] <= 0;
m[314] <= 0;
m[315] <= 0;
m[316] <= 0;
m[317] <= 0;
m[318] <= 0;
m[319] <= 0;
m[320] <= 0;
m[321] <= 0;
m[322] <= 0;
m[323] <= 0;
m[324] <= 0;
m[325] <= 0;
m[326] <= 0;
m[327] <= 0;
m[328] <= 0;
m[329] <= 0;
m[330] <= 0;
m[331] <= 0;
m[332] <= 0;
m[333] <= 0;
m[334] <= 0;
m[335] <= 0;
m[336] <= 0;
m[337] <= 0;
m[338] <= 0;
m[339] <= 0;
m[340] <= 0;
m[341] <= 0;
m[342] <= 0;
m[343] <= 0;
m[344] <= 0;
m[345] <= 0;
m[346] <= 0;
m[347] <= 0;
m[348] <= 0;
m[349] <= 0;
m[350] <= 0;
m[351] <= 0;
m[352] <= 0;
m[353] <= 0;
m[354] <= 0;
m[355] <= 0;
m[356] <= 0;
m[357] <= 0;
m[358] <= 0;
m[359] <= 0;
m[360] <= 0;
m[361] <= 0;
m[362] <= 0;
m[363] <= 0;
m[364] <= 0;
m[365] <= 0;
m[366] <= 0;
m[367] <= 0;
m[368] <= 0;
m[369] <= 0;
m[370] <= 0;
m[371] <= 0;
m[372] <= 0;
m[373] <= 0;
m[374] <= 0;
m[375] <= 0;
m[376] <= 0;
m[377] <= 0;
m[378] <= 0;
m[379] <= 0;
m[380] <= 0;
m[381] <= 0;
m[382] <= 0;
m[383] <= 0;
m[384] <= 0;
m[385] <= 0;
m[386] <= 0;
m[387] <= 0;
m[388] <= 0;
m[389] <= 0;
m[390] <= 0;
m[391] <= 0;
m[392] <= 0;
m[393] <= 0;
m[394] <= 0;
m[395] <= 0;
m[396] <= 0;
m[397] <= 0;
m[398] <= 0;
m[399] <= 0;
m[400] <= 0;
m[401] <= 0;
m[402] <= 0;
m[403] <= 0;
m[404] <= 0;
m[405] <= 0;
m[406] <= 0;
m[407] <= 0;
m[408] <= 0;
m[409] <= 0;
m[410] <= 0;
m[411] <= 0;
m[412] <= 0;
m[413] <= 0;
m[414] <= 0;
m[415] <= 0;
m[416] <= 0;
m[417] <= 0;
m[418] <= 0;
m[419] <= 0;
m[420] <= 0;
m[421] <= 0;
m[422] <= 0;
m[423] <= 0;
m[424] <= 0;
m[425] <= 0;
m[426] <= 0;
m[427] <= 0;
m[428] <= 0;
m[429] <= 0;
m[430] <= 0;
m[431] <= 0;
m[432] <= 0;
m[433] <= 0;
m[434] <= 0;
m[435] <= 0;
m[436] <= 0;
m[437] <= 0;
m[438] <= 0;
m[439] <= 0;
m[440] <= 0;
m[441] <= 0;
m[442] <= 0;
m[443] <= 0;
m[444] <= 0;
m[445] <= 0;
m[446] <= 0;
m[447] <= 0;
m[448] <= 0;
m[449] <= 0;
m[450] <= 0;
m[451] <= 0;
m[452] <= 0;
m[453] <= 0;
m[454] <= 0;
m[455] <= 0;
m[456] <= 0;
m[457] <= 0;
m[458] <= 0;
m[459] <= 0;
m[460] <= 0;
m[461] <= 0;
m[462] <= 0;
m[463] <= 0;
m[464] <= 0;
m[465] <= 0;
m[466] <= 0;
m[467] <= 0;
m[468] <= 0;
m[469] <= 0;
m[470] <= 0;
m[471] <= 0;
m[472] <= 0;
m[473] <= 0;
m[474] <= 0;
m[475] <= 0;
m[476] <= 0;
m[477] <= 0;
m[478] <= 0;
m[479] <= 0;
m[480] <= 0;
m[481] <= 0;
m[482] <= 0;
m[483] <= 0;
m[484] <= 0;
m[485] <= 0;
m[486] <= 0;
m[487] <= 0;
m[488] <= 0;
m[489] <= 0;
m[490] <= 0;
m[491] <= 0;
m[492] <= 0;
m[493] <= 0;
m[494] <= 0;
m[495] <= 0;
m[496] <= 0;
m[497] <= 0;
m[498] <= 0;
m[499] <= 0;
m[500] <= 0;
m[501] <= 0;
m[502] <= 0;
m[503] <= 0;
m[504] <= 0;
m[505] <= 0;
m[506] <= 0;
m[507] <= 0;
m[508] <= 0;
m[509] <= 0;
m[510] <= 0;
m[511] <= 0;
m[512] <= 0;
m[513] <= 0;
m[514] <= 0;
m[515] <= 0;
m[516] <= 0;
m[517] <= 0;
m[518] <= 0;
m[519] <= 0;
m[520] <= 0;
m[521] <= 0;
m[522] <= 0;
m[523] <= 0;
m[524] <= 0;
m[525] <= 0;
m[526] <= 0;
m[527] <= 0;
m[528] <= 0;
m[529] <= 0;
m[530] <= 0;
m[531] <= 0;
m[532] <= 0;
m[533] <= 0;
m[534] <= 0;
m[535] <= 0;
m[536] <= 0;
m[537] <= 0;
m[538] <= 0;
m[539] <= 0;
m[540] <= 0;
m[541] <= 0;
m[542] <= 0;
m[543] <= 0;
m[544] <= 0;
m[545] <= 0;
m[546] <= 0;
m[547] <= 0;
m[548] <= 0;
m[549] <= 0;
m[550] <= 0;
m[551] <= 0;
m[552] <= 0;
m[553] <= 0;
m[554] <= 0;
m[555] <= 0;
m[556] <= 0;
m[557] <= 0;
m[558] <= 0;
m[559] <= 0;
m[560] <= 0;
m[561] <= 0;
m[562] <= 0;
m[563] <= 0;
m[564] <= 0;
m[565] <= 0;
m[566] <= 0;
m[567] <= 0;
m[568] <= 0;
m[569] <= 0;
m[570] <= 0;
m[571] <= 0;
m[572] <= 0;
m[573] <= 0;
m[574] <= 0;
m[575] <= 0;
m[576] <= 0;
m[577] <= 0;
m[578] <= 0;
m[579] <= 0;
m[580] <= 0;
m[581] <= 0;
m[582] <= 0;
m[583] <= 0;
m[584] <= 0;
m[585] <= 0;
m[586] <= 0;
m[587] <= 0;
m[588] <= 0;
m[589] <= 0;
m[590] <= 0;
m[591] <= 0;
m[592] <= 0;
m[593] <= 0;
m[594] <= 0;
m[595] <= 0;
m[596] <= 0;
m[597] <= 0;
m[598] <= 0;
m[599] <= 0;
m[600] <= 0;
m[601] <= 0;
m[602] <= 0;
m[603] <= 0;
m[604] <= 0;
m[605] <= 0;
m[606] <= 0;
m[607] <= 0;
m[608] <= 0;
m[609] <= 0;
m[610] <= 0;
m[611] <= 0;
m[612] <= 0;
m[613] <= 0;
m[614] <= 0;
m[615] <= 0;
m[616] <= 0;
m[617] <= 0;
m[618] <= 0;
m[619] <= 0;
m[620] <= 0;
m[621] <= 0;
m[622] <= 0;
m[623] <= 0;
m[624] <= 0;
m[625] <= 0;
m[626] <= 0;
m[627] <= 0;
m[628] <= 0;
m[629] <= 0;
m[630] <= 0;
m[631] <= 0;
m[632] <= 0;
m[633] <= 0;
m[634] <= 0;
m[635] <= 0;
m[636] <= 0;
m[637] <= 0;
m[638] <= 0;
m[639] <= 0;
m[640] <= 0;
m[641] <= 0;
m[642] <= 0;
m[643] <= 0;
m[644] <= 0;
m[645] <= 0;
m[646] <= 0;
m[647] <= 0;
m[648] <= 0;
m[649] <= 0;
m[650] <= 0;
m[651] <= 0;
m[652] <= 0;
m[653] <= 0;
m[654] <= 0;
m[655] <= 0;
m[656] <= 0;
m[657] <= 0;
m[658] <= 0;
m[659] <= 0;
m[660] <= 0;
m[661] <= 0;
m[662] <= 0;
m[663] <= 0;
m[664] <= 0;
m[665] <= 0;
m[666] <= 0;
m[667] <= 0;
m[668] <= 0;
m[669] <= 0;
m[670] <= 0;
m[671] <= 0;
m[672] <= 0;
m[673] <= 0;
m[674] <= 0;
m[675] <= 0;
m[676] <= 0;
m[677] <= 0;
m[678] <= 0;
m[679] <= 0;
m[680] <= 0;
m[681] <= 0;
m[682] <= 0;
m[683] <= 0;
m[684] <= 0;
m[685] <= 0;
m[686] <= 0;
m[687] <= 0;
m[688] <= 0;
m[689] <= 0;
m[690] <= 0;
m[691] <= 0;
m[692] <= 0;
m[693] <= 0;
m[694] <= 0;
m[695] <= 0;
m[696] <= 0;
m[697] <= 0;
m[698] <= 0;
m[699] <= 0;
m[700] <= 0;
m[701] <= 0;
m[702] <= 0;
m[703] <= 0;
m[704] <= 0;
m[705] <= 0;
m[706] <= 0;
m[707] <= 0;
m[708] <= 0;
m[709] <= 0;
m[710] <= 0;
m[711] <= 0;
m[712] <= 0;
m[713] <= 0;
m[714] <= 0;
m[715] <= 0;
m[716] <= 0;
m[717] <= 0;
m[718] <= 0;
m[719] <= 0;
m[720] <= 0;
m[721] <= 0;
m[722] <= 0;
m[723] <= 0;
m[724] <= 0;
m[725] <= 0;
m[726] <= 0;
m[727] <= 0;
m[728] <= 0;
m[729] <= 0;
m[730] <= 0;
m[731] <= 0;
m[732] <= 0;
m[733] <= 0;
m[734] <= 0;
m[735] <= 0;
m[736] <= 0;
m[737] <= 0;
m[738] <= 0;
m[739] <= 0;
m[740] <= 0;
m[741] <= 0;
m[742] <= 0;
m[743] <= 0;
m[744] <= 0;
m[745] <= 0;
m[746] <= 0;
m[747] <= 0;
m[748] <= 0;
m[749] <= 0;
m[750] <= 0;
m[751] <= 0;
m[752] <= 0;
m[753] <= 0;
m[754] <= 0;
m[755] <= 0;
m[756] <= 0;
m[757] <= 0;
m[758] <= 0;
m[759] <= 0;
m[760] <= 0;
m[761] <= 0;
m[762] <= 0;
m[763] <= 0;
m[764] <= 0;
m[765] <= 0;
m[766] <= 0;
m[767] <= 0;
m[768] <= 0;
m[769] <= 0;
m[770] <= 0;
m[771] <= 0;
m[772] <= 0;
m[773] <= 0;
m[774] <= 0;
m[775] <= 0;
m[776] <= 0;
m[777] <= 0;
m[778] <= 0;
m[779] <= 0;
m[780] <= 0;
m[781] <= 0;
m[782] <= 0;
m[783] <= 0;
m[784] <= 0;
m[785] <= 0;
m[786] <= 0;
m[787] <= 0;
m[788] <= 0;
m[789] <= 0;
m[790] <= 0;
m[791] <= 0;
m[792] <= 0;
m[793] <= 0;
m[794] <= 0;
m[795] <= 0;
m[796] <= 0;
m[797] <= 0;
m[798] <= 0;
m[799] <= 0;
m[800] <= 0;
m[801] <= 0;
m[802] <= 0;
m[803] <= 0;
m[804] <= 0;
m[805] <= 0;
m[806] <= 0;
m[807] <= 0;
m[808] <= 0;
m[809] <= 0;
m[810] <= 0;
m[811] <= 0;
m[812] <= 0;
m[813] <= 0;
m[814] <= 0;
m[815] <= 0;
m[816] <= 0;
m[817] <= 0;
m[818] <= 0;
m[819] <= 0;
m[820] <= 0;
m[821] <= 0;
m[822] <= 0;
m[823] <= 0;
m[824] <= 0;
m[825] <= 0;
m[826] <= 0;
m[827] <= 0;
m[828] <= 0;
m[829] <= 0;
m[830] <= 0;
m[831] <= 0;
m[832] <= 0;
m[833] <= 0;
m[834] <= 0;
m[835] <= 0;
m[836] <= 0;
m[837] <= 0;
m[838] <= 0;
m[839] <= 0;
m[840] <= 0;
m[841] <= 0;
m[842] <= 0;
m[843] <= 0;
m[844] <= 0;
m[845] <= 0;
m[846] <= 0;
m[847] <= 0;
m[848] <= 0;
m[849] <= 0;
m[850] <= 0;
m[851] <= 0;
m[852] <= 0;
m[853] <= 0;
m[854] <= 0;
m[855] <= 0;
m[856] <= 0;
m[857] <= 0;
m[858] <= 0;
m[859] <= 0;
m[860] <= 0;
m[861] <= 0;
m[862] <= 0;
m[863] <= 0;
m[864] <= 0;
m[865] <= 0;
m[866] <= 0;
m[867] <= 0;
m[868] <= 0;
m[869] <= 0;
m[870] <= 0;
m[871] <= 0;
m[872] <= 0;
m[873] <= 0;
m[874] <= 0;
m[875] <= 0;
m[876] <= 0;
m[877] <= 0;
m[878] <= 0;
m[879] <= 0;
m[880] <= 0;
m[881] <= 0;
m[882] <= 0;
m[883] <= 0;
m[884] <= 0;
m[885] <= 0;
m[886] <= 0;
m[887] <= 0;
m[888] <= 0;
m[889] <= 0;
m[890] <= 0;
m[891] <= 0;
m[892] <= 0;
m[893] <= 0;
m[894] <= 0;
m[895] <= 0;
m[896] <= 0;
m[897] <= 0;
m[898] <= 0;
m[899] <= 0;
m[900] <= 0;
m[901] <= 0;
m[902] <= 0;
m[903] <= 0;
m[904] <= 0;
m[905] <= 0;
m[906] <= 0;
m[907] <= 0;
m[908] <= 0;
m[909] <= 0;
m[910] <= 0;
m[911] <= 0;
m[912] <= 0;
m[913] <= 0;
m[914] <= 0;
m[915] <= 0;
m[916] <= 0;
m[917] <= 0;
m[918] <= 0;
m[919] <= 0;
m[920] <= 0;
m[921] <= 0;
m[922] <= 0;
m[923] <= 0;
m[924] <= 0;
m[925] <= 0;
m[926] <= 0;
m[927] <= 0;
m[928] <= 0;
m[929] <= 0;
m[930] <= 0;
m[931] <= 0;
m[932] <= 0;
m[933] <= 0;
m[934] <= 0;
m[935] <= 0;
m[936] <= 0;
m[937] <= 0;
m[938] <= 0;
m[939] <= 0;
m[940] <= 0;
m[941] <= 0;
m[942] <= 0;
m[943] <= 0;
m[944] <= 0;
m[945] <= 0;
m[946] <= 0;
m[947] <= 0;
m[948] <= 0;
m[949] <= 0;
m[950] <= 0;
m[951] <= 0;
m[952] <= 0;
m[953] <= 0;
m[954] <= 0;
m[955] <= 0;
m[956] <= 0;
m[957] <= 0;
m[958] <= 0;
m[959] <= 0;
m[960] <= 0;
m[961] <= 0;
m[962] <= 0;
m[963] <= 0;
m[964] <= 0;
m[965] <= 0;
m[966] <= 0;
m[967] <= 0;
m[968] <= 0;
m[969] <= 0;
m[970] <= 0;
m[971] <= 0;
m[972] <= 0;
m[973] <= 0;
m[974] <= 0;
m[975] <= 0;
m[976] <= 0;
m[977] <= 0;
m[978] <= 0;
m[979] <= 0;
m[980] <= 0;
m[981] <= 0;
m[982] <= 0;
m[983] <= 0;
m[984] <= 0;
m[985] <= 0;
m[986] <= 0;
m[987] <= 0;
m[988] <= 0;
m[989] <= 0;
m[990] <= 0;
m[991] <= 0;
m[992] <= 0;
m[993] <= 0;
m[994] <= 0;
m[995] <= 0;
m[996] <= 0;
m[997] <= 0;
m[998] <= 0;
m[999] <= 0;
m[1000] <= 0;
m[1001] <= 0;
m[1002] <= 0;
m[1003] <= 0;
m[1004] <= 0;
m[1005] <= 0;
m[1006] <= 0;
m[1007] <= 0;
m[1008] <= 0;
m[1009] <= 0;
m[1010] <= 0;
m[1011] <= 0;
m[1012] <= 0;
m[1013] <= 0;
m[1014] <= 0;
m[1015] <= 0;
m[1016] <= 0;
m[1017] <= 0;
m[1018] <= 0;
m[1019] <= 0;
m[1020] <= 0;
m[1021] <= 0;
m[1022] <= 0;
m[1023] <= 0;
	end
end


endmodule
