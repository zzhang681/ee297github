
module img_ram_test (
	address,
	clock,
	data,
	wren,
	q
);

input	[9:0]  address;
	input	  clock;
	input	[7:0]  data;
	input	  wren;
	output	[7:0]  q;








endmodule
