// fp_mac.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module fp_mac (
		input  wire        clk,       // s1.clk
		input  wire			 clk_50,
		input  [127:0]		 data,
		input  wire [31:0] din,			//input(image)
		input  wire	[31:0] din_bias,
		input					 datavalid,
		input  wire        reset,     //   .reset
		input  wire        start,     //   .start
		input 	[9:0]		 i_addr_r,
		input  wire [127:0] interface_address,
		input  wire 			empty,
		output logic        ready,      //   .ready
		output reg [3:0] index_pred,
		output wire [31:0] result,     //   .result
		output wire [4:0] states,
		output wire next_in,
		output adone
		
);

enum bit[4:0] {
	IDLE,				//Stay Idle until Reader finished loading image into SRAM
	READ_IMG,		//not used
	OP_START,		//Send read request to FIFO, wait weight data
	READ,				//not used
	READ_DONE,		//not used
	OP,				//Perform multiplication & Accumulation for 1 group of weight data
	OP_DONE,			//Finish buffer state, store result into hidden SRAM
	BIAS_START,		//00111
	BIAS,				//01000
	BIAS_DONE,		//01001
	RELU_START,		//01010
	RELU,				//01011
	HO_READ_START,		//01100
	HO_OP_START,				//01101
	HO_OP,		//01110
	HO_OP1_DONE,
	HO_OP2,
	HO_OP_DONE,			//10000
	HO_BIAS_START,
	HO_BIAS,
	HO_BIAS1_DONE,
	HO_BIAS2,
	HO_BIAS_DONE,
	HO_RELU,
	OUT_BUFFER,
	OUT_COMPARE,
	ALL_DONE			//10001
} cs, ns;

assign count_ho_ob = count_ho;

//typedef union packed{
//logic [63:0][31:0] h;
//} hidden_reg;

assign states = cs;
//hidden_reg hidden;


logic [31:0] dataa_bias, datab_bias, result_bias;
logic start_bias;
logic [7:0] count_bias;

logic [5:0] count_ho;
logic [63:0] wdata_ho,rdata_ho;
logic [3:0] addr_w_ho,addr_r_ho;
logic write_ho, read_ho;
logic [127:0] weight_reg_ho;
logic highbit_ho;

parameter ADDR_W1 = 0;
parameter ADDR_W1_FIN = 200703;
parameter ADDR_BIAS1 = 200704;
parameter ADDR_BIAS1_FIN = 200959;
parameter ADDR_W2 = 200960;
parameter ADDR_W2_FIN = 203519;
parameter ADDR_BIAS2 = 203520;
parameter ADDR_BIAS2_FIN = 203559;

parameter COUNT_ACC_CYCLE = 5;



logic [31:0] dataa1, datab1, result_mul1;
logic [31:0] dataa2, datab2, result_mul2;
logic [31:0] dataa3, datab3, result_mul3;
logic [31:0] dataa4, datab4, result_mul4;

logic [31:0] dataa1_add, datab1_add;
logic [31:0] dataa2_add, datab2_add;
logic [31:0] dataa3_add, datab3_add;
logic [31:0] dataa4_add, datab4_add;
logic [31:0] result_add1, result_add2, result_add3, result_add4;
logic [127:0] result_add_reg;

logic done_mul1;
logic done_mul2;
logic done_mul3;
logic done_mul4;
logic done_flag1, done_flag2, done_flag3, done_flag4;

logic [31:0] x0,x1,x2,x3;//, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15;
logic [31:0] r0,r1,r2,r3;//, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15;
logic [3:0] n0;//, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;
//logic [3:0] acc_en0, acc_en1, acc_en2, acc_en3, acc_en4, acc_en5, acc_en6, acc_en7, acc_en8, acc_en9, acc_en10, acc_en11, acc_en12, acc_en13, acc_en14, acc_en15;

//logic []

logic we, re;

//logic [2:0] n_mul, n_add;
logic clk_en, reset_req;
logic [3:0] address, address_next;		//address for hidden (0-63)
logic address_hidden_read;

logic [3:0] count_mul;

logic next_in_edge, done_re_level;
logic start_mul;
logic next_address_ready;
logic next_in_ho;
assign edge_det_READ = (cs == READ) ? 1:0;
assign adone = (cs == ALL_DONE) ? 1:0;
assign next_in = (address == 15) & (cs == OP_DONE);
assign next_in_ho = (address_ho == 4) & (cs == HO_OP_DONE || cs == HO_OP1_DONE);

logic [127:0] wdata_hidden, rdata_hidden;
logic wren_hidden;
logic [4:0] address_hidden;
logic [3:0] count;
logic [31:0] count_num_mul;


logic [3:0] address_ho, address_ho_next;		//hidden - out, 0-4


logic [5:0] address_out;
logic [63:0] wdata_out, rdata_out;
logic wren_out;


//assign reset_req = !reset;//(cs == IDLE) ? 1:0;

/*
assign dataa_fp = 32'h3e99999a;	//0.3
assign datab_fp = 32'h3ecccccd;	//0.4		//expect multiply result 0.12 3df5c28f
*/


parameter n_mul = 3'b100;
parameter n_add = 3'b101;
//multiply: 100
//add: 101

assign clk_en = 1'b1;

always @(*) begin
	ready = 0;
	begin
		case(cs)
			IDLE: ready = 0;
			OP_START: begin 
				if(count == 0) ready = 1;
				else ready = 0;
			end
			OP: begin 
					ready = 0; 
			end
			BIAS_START: begin
				if(count == 0) ready = 1;
				else ready = 0;
			end
			HO_OP_START: begin 
				if(count == 0) ready = 1;
				else ready = 0;
			end
			HO_OP: ready = 0;
			HO_BIAS_START: begin
				if(count == 0) ready = 1;
				else ready = 0;
			end
			//OP_DONE: ready = 1;
			default: ready = 0;
		endcase
	end
end
	

//count 5 cycles and store the result///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//add a sram to store hidden
always @(posedge clk) begin
	if(reset) count <= 0;
	else begin
		if(cs == OP_START) begin
			case(count)
				0: if(!empty) count <= count + 1;
				1: count <= 0;
			endcase
		end else if(cs == OP) begin
		case(count)
			0: begin
				if(done_mul1) count <= count + 1;
				else count <= 0;
			end
			COUNT_ACC_CYCLE: begin
				count <= 0;
			end
			default: count <= count + 1;
		endcase
		end else if(cs == BIAS_START) begin
			case(count)
				0: if(!empty) count <= count + 1;
				1: count <= 0;
			endcase
		end else if(cs == BIAS) begin
		case(count)
			0: begin
				count <= count + 1;
			end
			COUNT_ACC_CYCLE: begin
				count <= 0;
			end
			default: count <= count + 1;
		endcase
		end
		else if(cs == RELU) begin
			case(count)
				0: begin
					count <= count + 1;
				end
				2: count <= 0;
				default: count <= count + 1;
			endcase
		end
		else if(cs == HO_OP_START) begin
			case(count)
				0: if(!empty) count <= count + 1;
				1: count <= 0;
			endcase
		end else if(cs == HO_OP) begin
		case(count)
			0: begin
				if(done_mul1) count <= count + 1;
				else count <= 0;
			end
			COUNT_ACC_CYCLE: begin
				count <= 0;
			end
			default: count <= count + 1;
		endcase
		end else if(cs == HO_OP2) begin
		case(count)
			0: begin
				if(done_mul1) count <= count + 1;
				else count <= 0;
			end
			COUNT_ACC_CYCLE: begin
				count <= 0;
			end
			default: count <= count + 1;
		endcase
		end else if(cs == HO_BIAS_START) begin
			case(count)
				0: if(!empty) count <= count + 1;
				1: count <= 0;
			endcase
		end else if(cs == HO_BIAS) begin
		case(count)
			0: begin
				count <= count + 1;
			end
			COUNT_ACC_CYCLE: begin
				count <= 0;
			end
			default: count <= count + 1;
		endcase
		end else if(cs == HO_BIAS2) begin
		case(count)
			0: begin
				count <= count + 1;
			end
			COUNT_ACC_CYCLE: begin
				count <= 0;
			end
			default: count <= count + 1;
		endcase
		end
		else if(cs == HO_RELU) begin
			case(count)
				0: begin
					count <= count + 1;
				end
				2: count <= 0;
				default: count <= count + 1;
			endcase
		end 
		else if(cs == OUT_COMPARE) begin
			case(count)
				0: begin
					count <= count + 1;
				end
				3: count <= 0;
				default: count <= count + 1;
			endcase
		end 
	end
end


//count_bias

/*
1. start -> 9 cycle -> done -> wait start   (Finished)
2. make sure read correctly    (Finished?)
3. 1 IP start -> wait done			(Finished)
4. make sure result correct with mul & add with simple inputs	(Finished)
5. ****try some new inputs read from SDRAM****                  (Finished)
0 -> 0.1   16 -> 0.2    32 -> 0.3     48 -> 0.4    64 -> 0.5
3DCCCCCD   3E4CCCCD 32  3E99999A 48   3ECCCCCD     3F000000
in: 0.5       16   32  48   64
result: 0.05+0.1+0.15+0.2+0.25=0.75 (3F400000)
0.95 (0.75) (+0.2)
0.65 (0.5)  (+0.15)
0.4  (0.3)  (+0.1)  (0.05+0.1+0.15+0.1)
0.2  (0.15) (+0.05) (0.05+0.1+0.05)
6. PROBLEM: hidden: no reset problem? (Finished, final address may different)
7. Check m2-m4 stability   (Finished)
8. Add states to update input
	problem: unstable
	single input: finished
	different inputs
		something wrong with the input change (Finished)
9. how to input image?           (Finished)
	address 204000 - 204783
10. address of image does not increase
10.5. add bias
11. add ReLU
*/

//ns
always_comb begin
	ns = cs;
	case(cs)
		IDLE: begin
			if(start) ns = OP_START;
			else ns = IDLE;
		end
		
		OP_START: begin
			if(count == 1) ns = OP;
			else ns = OP_START;
		end
		
		OP: begin
			if(done_flag1 && done_flag2 && done_flag3 &&done_flag4 && count == COUNT_ACC_CYCLE) begin
				ns = OP_DONE;
			end else ns = OP;
		end
		
		OP_DONE: begin 
			if(interface_address >= ADDR_BIAS1 && empty) ns = BIAS_START;
			else ns = OP_START;
		end
		
		BIAS_START: begin
			if(count == 1) ns = BIAS;
			else ns = BIAS_START;
		end
		
		BIAS: begin
			if(count == COUNT_ACC_CYCLE) ns = BIAS_DONE;
			else ns = BIAS;
		end
		
		BIAS_DONE: begin
			if(interface_address >= ADDR_W2 && empty) ns = RELU;
			else ns = BIAS_START;
		end
		
		RELU: begin
			if(address == 15 && count == 2) ns = HO_OP_START;
			else ns = RELU;
		end
		HO_OP_START: begin
			if(count == 1) ns = HO_OP;
			else ns = HO_OP_START;
		end
		
		HO_OP: begin
			if(done_flag1 && done_flag2 && count == COUNT_ACC_CYCLE) begin
				ns = HO_OP1_DONE;
			end else ns = HO_OP;
		end
		HO_OP1_DONE: begin
			if(count_ho >= 63 && address_ho >= 4) ns = HO_BIAS_START;
			else ns = HO_OP2;
		end
		HO_OP2: begin
			if(done_flag1 && count == COUNT_ACC_CYCLE) begin
				ns = HO_OP_DONE;
			end else ns = HO_OP2;
		end
		HO_OP_DONE: begin
			if(count_ho >= 63 && address_ho >= 4) ns = HO_BIAS_START;
			else ns = HO_OP_START;
		end
		HO_BIAS_START: begin
			if(count == 1) ns = HO_BIAS;
			else ns = HO_BIAS_START;
		end
		HO_BIAS: begin
			if(count == COUNT_ACC_CYCLE) ns = HO_BIAS1_DONE;
			else ns = HO_BIAS;
		end
		HO_BIAS1_DONE: begin
			if(empty) ns = HO_RELU;
			else ns = HO_BIAS2;
		end
		HO_BIAS2: begin
			if(count == COUNT_ACC_CYCLE) ns = HO_BIAS_DONE;
			else ns = HO_BIAS2;
		end
		HO_BIAS_DONE: begin
			if(empty) ns = HO_RELU;
			else ns = HO_BIAS_START;
		end
		HO_RELU: begin
			if(address_out == 4 && count == 2) ns = OUT_BUFFER;
			else ns = HO_RELU;
		end
		OUT_BUFFER: ns = OUT_COMPARE;
		OUT_COMPARE: begin
			if(address_out == 4 && count == 3) ns = ALL_DONE;
			else ns = OUT_COMPARE;
		end
		ALL_DONE: ns = ALL_DONE;
		
	endcase
end

// ----------------------- CONTROL SIGNALS ------------------------- //
//start_mul
/*
always @(posedge clk) begin
	if(reset) start_mul <= 0;
	else if(datavalid && done) start_mul <= 1;
end
*/


always @(posedge clk) begin
	if(reset) start_mul <= 0;
	else if(cs == OP_START && ns == OP) start_mul <= 1;
	else if(cs == HO_OP_START && ns == HO_OP)start_mul <= 1;
	else if(cs == HO_OP1_DONE && ns == HO_OP2) start_mul <= 1;
	else start_mul <= 0;
end

//count_mul
always @(posedge clk) begin
	if(reset) count_mul <= 0;
	else begin
	if(cs == OP) begin
		case(count_mul)
			0: begin
				if(start_mul) count_mul <= count_mul + 1;
				else count_mul <= 0;
			end
			4: count_mul <= 0;
			default: count_mul <= count_mul + 1;
		endcase
	end else if(cs == HO_OP || cs == HO_OP2) begin
		case(count_mul)
			0: begin
				if(start_mul) count_mul <= count_mul + 1;
				else count_mul <= 0;
			end
			4: count_mul <= 0;
			default: count_mul <= count_mul + 1;
		endcase
	end
	end
end

always @(*) begin
	done_mul1 = 0;
	done_mul2 = 0;
	if(cs == OP) begin
		if(count_mul == 3) begin
			done_mul1 = 1;
			done_mul2 = 1;
		end
	end else if(cs == HO_OP || cs == HO_OP2) begin
		if(count_mul == 4) begin
			done_mul1 = 1;
			done_mul2 = 1;
		end
	end
end
assign done_mul3 = count_mul == 3 ? 1:0;
assign done_mul4 = count_mul == 3 ? 1:0;


//address
always_ff @(posedge clk) begin
	if(reset) begin 
		address <= 0;
		address_ho <= 0;
	end else begin
		address <= address_next;
		address_ho <= address_ho_next;
	end
end

//address_next
always_comb begin
	address_next = address;
	address_ho_next = address_ho;
	case(cs)
		IDLE: begin
			address_next = 0;
			address_ho_next = 0;
		end
		OP_DONE: begin
			if(address<15) address_next = address + 1;
			else address_next = 0;
		end
		
		BIAS_DONE: begin
			if(address<15) address_next = address + 1;
			else address_next = 0;
		end
		
		RELU: begin
			if(count == 2) address_next = address + 1;
		end
		
		HO_OP_DONE: begin 
			if(address_ho < 4) address_ho_next = address_ho + 1;
			else address_ho_next = 0;
			
		end
		
		HO_OP1_DONE: begin 
			if(address_ho < 4) address_ho_next = address_ho + 1;
			else address_ho_next = 0;
		end
		
		HO_BIAS1_DONE: begin
			if(address_ho < 4) address_ho_next = address_ho + 1;
			else address_ho_next = 0;
		end
		
		HO_BIAS_DONE: begin
			if(address_ho < 4) address_ho_next = address_ho + 1;
			else address_ho_next = 0;
		end
		
		HO_RELU: begin
			if(count == 2) begin 
				if(address < 4) address_ho_next = address_ho + 1;
				else address_ho_next = 0;
			end
		end
		OUT_BUFFER: address_ho_next = 0;
		
		OUT_COMPARE: begin
			if(count == 3) address_ho_next = address_ho + 1;
		end
		
	endcase
end

assign address_hidden_read = 0;

always @(posedge clk) begin
	if(reset) begin
		done_flag1 <= 0;
		done_flag2 <= 0;
		done_flag3 <= 0;
		done_flag4 <= 0;
	end else begin
		if(done_mul1) done_flag1 <= 1;
		if(done_mul2) done_flag2 <= 1;
		if(done_mul3) done_flag3 <= 1;
		if(done_mul4) done_flag4 <= 1;
		if(cs != ns/*cs == OP_DONE*/) begin
			done_flag1 <= 0;
			done_flag2 <= 0;
			done_flag3 <= 0;
			done_flag4 <= 0;
		end
	end
end



//n = Boolean port which signals the beginning of a 
//new data set to be accumulated. This should go high 
//together with the first element in the new data set 
//and should go low the next cycle. The data sets may be 
//of variable length and a new data set may be started 
//at any time. The accumulation result for an input 
//is available after the reported latency. 


//count_ho
always @(posedge clk) begin
	if(reset) count_ho <= 0;
	else begin
		if(next_in_ho) begin
			count_ho <= count_ho + 1;
		end
	end
end

//count_num_mul
always @(posedge clk) begin
	if(reset) count_num_mul <= 0;
	else begin
		if(cs == HO_OP1_DONE || cs == HO_OP_DONE) begin
			count_num_mul <= count_num_mul + 2;
		end
	end
end



// ----------------------------------------------------------------- //


// ------------------------- DATA SIGNALS -------------------------- //////////////////////////////////////////////////////

logic [31:0] dataa_comp, datab_comp;
logic [31:0] reg_comp;
logic [3:0] index_comp;
logic [0:0] q_comp;
//logic [3:0] index_pred;

//assign index_pred1 = index_pred;

//dataa_comp, datab_comp
always @(*) begin
	dataa_comp = 0;
	datab_comp = 0;
	case(cs)
		OUT_COMPARE: begin
			case(count)
				2: begin
					dataa_comp = rdata_out[31:0];
					datab_comp = reg_comp;
				end
				3: begin
					dataa_comp = rdata_out[63:32];
					datab_comp = reg_comp;
				end
				default: begin
					dataa_comp = 0;
					datab_comp = 0;
				end
			endcase
		end
	endcase
end

always @(*) begin
	index_comp = 0;
	case(cs)
		OUT_COMPARE: begin
			if(count == 2) index_comp = address_out * 2;
			else if(count == 3) index_comp = address_out * 2 + 1;
		end
	endcase
end

always @(posedge clk) begin
	if(reset) begin
		reg_comp <= 0;
		index_pred <= 0;
	end else begin
		case(cs)
			OUT_COMPARE: begin
				case(count)
					2: begin
						//index_comp <= index_comp + 1;
						if(q_comp) begin
							reg_comp <= dataa_comp;
							index_pred <= index_comp;
						end else begin
							reg_comp <= datab_comp;
						end
					end
					3: begin
						//index_comp <= index_comp + 1;
						if(q_comp) begin
							reg_comp <= dataa_comp;
							index_pred <= index_comp;
						end else begin
							reg_comp <= datab_comp;
						end
					end
					default: begin
						//index_comp <= index_comp;
						index_pred <= index_pred;
						reg_comp <= reg_comp;
					end
				endcase
			end
			default: begin
				//index_comp <= index_comp;
				index_pred <= index_pred;
				reg_comp <= reg_comp;
			end
		endcase
	end
end





//assign start_add = done_mul1;
always @(*) begin
	start_add = 0;
	case(cs)
		OP: start_add = done_mul1;
		BIAS: begin
			if(count == 0) start_add = 1;
		end
		HO_OP: start_add = done_mul1;
		HO_OP2: start_add = done_mul1;
		HO_BIAS: begin
			if(count == 0) start_add = 1;
		end
		HO_BIAS2: begin
			if(count == 0) start_add = 1;
		end
	endcase
end


always @(*) begin
	dataa1_add = 0;
	datab1_add = 0;
	dataa2_add = 0;
	datab2_add = 0;
	dataa3_add = 0;
	datab3_add = 0;
	dataa4_add = 0;
	datab4_add = 0;
	case(cs)
		OP: begin
			//if(start_add) begin
				if(i_addr_r < 1) begin
					dataa1_add = 0;
					datab1_add = result_mul1;
					dataa2_add = 0;
					datab2_add = result_mul2;
					dataa3_add = 0;
					datab3_add = result_mul3;
					dataa4_add = 0;
					datab4_add = result_mul4;
				end else begin 
					dataa1_add = rdata_hidden[31:0];
					datab1_add = result_mul1;
					dataa2_add = rdata_hidden[63:32];
					datab2_add = result_mul2;
					dataa3_add = rdata_hidden[95:64];
					datab3_add = result_mul3;
					dataa4_add = rdata_hidden[127:96];
					datab4_add = result_mul4;
				end
			//end
		end
		BIAS: begin
			if(start_add) begin
				dataa1_add = rdata_hidden[31:0];
				datab1_add = data[31:0];
				dataa2_add = rdata_hidden[63:32];
				datab2_add = data[63:32];
				dataa3_add = rdata_hidden[95:64];
				datab3_add = data[95:64];
				dataa4_add = rdata_hidden[127:96];
				datab4_add = data[127:96];
			end
		end
		HO_OP: begin
			//if(start_add) begin
				if(count_ho < 1) begin
					dataa1_add = 0;
					datab1_add = result_mul1;
					dataa2_add = 0;
					datab2_add = result_mul2;
				end else begin 
					dataa1_add = rdata_out[31:0];
					datab1_add = result_mul1;
					dataa2_add = rdata_out[63:32];
					datab2_add = result_mul2;
				end
			//end
		end
		HO_OP2: begin
			//if(start_add) begin
				if(count_ho < 1) begin
					dataa1_add = 0;
					datab1_add = result_mul1;
					dataa2_add = 0;
					datab2_add = result_mul2;
				end else begin 
					dataa1_add = rdata_out[31:0];
					datab1_add = result_mul1;
					dataa2_add = rdata_out[63:32];
					datab2_add = result_mul2;
				end
			//end
		end
		HO_BIAS: begin
			if(start_add) begin
				dataa1_add = rdata_out[31:0];
				datab1_add = data[31:0];
				dataa2_add = rdata_out[63:32];
				datab2_add = data[63:32];
			end
		end
		HO_BIAS2: begin
			if(start_add) begin
				dataa1_add = rdata_out[31:0];
				datab1_add = data[95:64];
				dataa2_add = rdata_out[63:32];
				datab2_add = data[127:96];
			end
		end
	endcase
end

//result_add_reg
always @(posedge clk) begin
	if(reset) result_add_reg <= 0;
	else begin
		case(cs)
			OP: begin
				if(done_add1) result_add_reg[31:0] <= result_add1;
				if(done_add2) result_add_reg[63:32] <= result_add2;
				if(done_add3) result_add_reg[95:64] <= result_add3;
				if(done_add4) result_add_reg[127:96] <= result_add4;
			end
			OP_DONE: begin
				result_add_reg <= 0;
			end
		endcase
	end
end

logic [127:0] relu_temp;
always @(*) begin
	relu_temp = 0;
	if(cs == RELU) begin 
		relu_temp[127:96] = (rdata_hidden[127] == 1) ? 0 : rdata_hidden[127:96];
		relu_temp[95:64] = (rdata_hidden[95] == 1) ? 0 : rdata_hidden[95:64];
		relu_temp[63:32] = (rdata_hidden[63] == 1) ? 0 : rdata_hidden[63:32];
		relu_temp[31:0] = (rdata_hidden[31] == 1) ? 0 : rdata_hidden[31:0];
	end
end

logic [63:0] relu_temp_ho;
always @(*) begin
	relu_temp_ho = 0;
	if(cs == HO_RELU) begin 
		relu_temp_ho[63:32] = (rdata_out[63] == 1) ? 0 : rdata_out[63:32];
		relu_temp_ho[31:0] = (rdata_out[31] == 1) ? 0 : rdata_out[31:0];
	end
end

//hidden ram
always @(*) begin
	wdata_hidden = 0;
	wren_hidden = 0;
	address_hidden = 0;
	case(cs)
		OP_START: begin
			wren_hidden = 0;
			address_hidden = address;
		end
		OP: begin
			address_hidden = address;
		end
		OP_DONE: begin
			wren_hidden = 1;
			address_hidden = address;
			wdata_hidden = result_add_reg;//{r3,r2,r1,r0};
		end
		BIAS_START: begin
			wren_hidden = 0;
			address_hidden = address;
		end
		BIAS: begin
			address_hidden = address;
		end
		BIAS_DONE: begin
			wren_hidden = 1;
			address_hidden = address;
			wdata_hidden = rdata_hidden;
		end
		RELU: begin 
			address_hidden = address;
			if(count == 2) begin
				wren_hidden = 1;
				wdata_hidden = relu_temp;
			end
		end
		HO_OP_START: address_hidden = count_ho / 4;
		HO_OP: address_hidden = count_ho / 4;
		HO_OP1_DONE: address_hidden = count_ho / 4;
		HO_OP2: address_hidden = count_ho / 4;
		HO_OP_DONE: address_hidden = count_ho / 4;
		ALL_DONE: address_hidden = 0;
	endcase
end

//output ram
//[5:0] address_out;
//[63:0] wdata_out, rdata_out;
//wren_out;
always @(*) begin
	address_out = 0;
	wdata_out = 0;
	wren_out = 0;
	case(cs)
		HO_OP_START: begin
			wren_out = 0;
			address_out = address_ho;
		end
		HO_OP: address_out = address_ho;
		
		HO_OP1_DONE: begin
			wren_out = 1;
			address_out = address_ho;
			wdata_out = {result_add2, result_add1};
		end
		HO_OP2: address_out = address_ho;
		HO_OP_DONE: begin
			wren_out = 1;
			address_out = address_ho;
			wdata_out = {result_add2, result_add1};
		end
		HO_BIAS_START: address_out = address_ho;
		HO_BIAS: begin
			address_out = address_ho;
		end
		HO_BIAS1_DONE: begin
			wren_out = 1;
			address_out = address_ho;
			wdata_out = rdata_out;
		end
		HO_BIAS2: begin
			address_out = address_ho;
		end
		HO_BIAS_DONE: begin
			wren_out = 1;
			address_out = address_ho;
			wdata_out = rdata_out;
		end
		HO_RELU: begin 
			address_out = address_ho;
			if(count == 2) begin
				wren_out = 1;
				wdata_out = relu_temp_ho;
			end
		end
		OUT_COMPARE: begin
			address_out = address_ho;
		end
	endcase
end



//x15;
always @(*) begin
	x0 = 0;
	x1 = 0;
	x2 = 0;
	x3 = 0;
	case(cs)
		OP_START: begin
			if(ns == OP) begin
				if(i_addr_r < 1) begin
					x0 = 0;
					x1 = 0;
					x2 = 0;
					x3 = 0;
				end else begin 
					x0 = rdata_hidden[31:0];
					x1 = rdata_hidden[63:32];
					x2 = rdata_hidden[95:64];
					x3 = rdata_hidden[127:96];
				end
			end
		end
		OP: begin
			if(done_mul1) x0 = result_mul1;
			if(done_mul2) x1 = result_mul2;
			if(done_mul3) x2 = result_mul3;
			if(done_mul4) x3 = result_mul4;
		end
		
	endcase
end
	

//dataa1 - 4. datab1 - 4
always @(*) begin
	dataa1 = 0;
	dataa2 = 0;
	dataa3 = din;
	dataa4 = din;
	datab1 = 0;
	datab2 = 0;
	datab3 = 0;
	datab4 = 0;
	case(cs)
		OP_START: begin
			dataa1 = din;
			dataa2 = din;
			datab1 = data[31:0];
			datab2 = data[63:32];
			datab3 = data[95:64];
			datab4 = data[127:96];
		end
		OP: begin
			dataa1 = din;
			dataa2 = din;
			datab1 = data[31:0];
			datab2 = data[63:32];
			datab3 = data[95:64];
			datab4 = data[127:96];
		end
		HO_OP: begin
			datab1 = weight_reg_ho[31:0];
			datab2 = weight_reg_ho[63:32];
			case(count_ho % 4)
				0: begin
					dataa1 = rdata_hidden[31:0];
					dataa2 = rdata_hidden[31:0];
				end
				1: begin
					dataa1 = rdata_hidden[63:32];
					dataa2 = rdata_hidden[63:32];
				end
				2: begin
					dataa1 = rdata_hidden[95:64];
					dataa2 = rdata_hidden[95:64];
				end
				3: begin
					dataa1 = rdata_hidden[127:96];
					dataa2 = rdata_hidden[127:96];
				end
			endcase
		end
		HO_OP2: begin
			datab1 = weight_reg_ho[95:64];
			datab2 = weight_reg_ho[127:96];
			case(count_ho % 4)
				0: begin
					dataa1 = rdata_hidden[31:0];
					dataa2 = rdata_hidden[31:0];
				end
				1: begin
					dataa1 = rdata_hidden[63:32];
					dataa2 = rdata_hidden[63:32];
				end
				2: begin
					dataa1 = rdata_hidden[95:64];
					dataa2 = rdata_hidden[95:64];
				end
				3: begin
					dataa1 = rdata_hidden[127:96];
					dataa2 = rdata_hidden[127:96];
				end
			endcase
		end
	endcase
end



//weight_reg_ho
always @(posedge clk) begin
	if(reset) weight_reg_ho <= 0;
	else begin
		if(datavalid && cs == HO_OP_START) weight_reg_ho <= data;
	end
end

//wdata_ho


//highbit_ho
always @(posedge clk) begin
	if(reset) highbit_ho <= 0;
	else begin
		if(cs == HO_OP) begin
			case(highbit_ho)
				0: begin
					if(done_mul1) highbit_ho <= 1;
				end
				1: begin
					if(done_mul1) highbit_ho <= 0;
				end
			endcase
		end
	end
end



// ----------------------------------------------------------------- //

// ------------------------- TEST SIGNALS -------------------------- //

logic [31:0] data_test;

always_ff @(posedge clk) begin
	if(reset) data_test <= 0;
	else begin
		data_test <= address;//r0[31:0];//rdata_ho[31:0];////i_addr_r;//datab1;//result_add1;//din;////result_add1;
	end
end

//result


always_ff @(posedge clk) begin
	if(reset) result <= 0;
	else begin
		result <= data_test;//hidden[0][31:0];//dataa1;//result_add1;//din;//hidden[0][31:0];//result_add1;
	end
end

logic [9:0] wf_count;

always_ff @(posedge clk) begin
	if(reset) wf_count <= 0;
	else begin
			if(next_in_edge) wf_count <= wf_count + 1;			//count how many ops in total
			else wf_count <= wf_count;
	end
end


//assign result = result_bias;//count_bias;//address;


// ----------------------------------------------------------------- //



//cs
always_ff @(posedge clk) begin
	if(reset) cs <= IDLE;
	else cs <= ns;
end

//4 muls

fptest fp1(
	.clk(clk),
	.areset(reset),
	.en(1'b1),
	.a(dataa1),
	.b(datab1),
	.q(result_mul1)
);

fptest fp2(
	.clk(clk),
	.areset(reset),
	.en(1'b1),
	.a(dataa2),
	.b(datab2),
	.q(result_mul2)
);

fptest fp3(
	.clk(clk),
	.areset(reset),
	.en(1'b1),
	.a(dataa3),
	.b(datab3),
	.q(result_mul3)
);

fptest fp4(
	.clk(clk),
	.areset(reset),
	.en(1'b1),
	.a(dataa4),
	.b(datab4),
	.q(result_mul4)
);

//muls



fpoint2_multi #(
		.arithmetic_present (1),
		.root_present       (1),
		.conversion_present (1)
	) nios_custom_instr_floating_point_2_multi_1 (
		.clk       (clk),       // s1.clk
		.clk_en    (clk_en),    //   .clk_en
		.dataa     (dataa1_add),     //   .dataa
		.datab     (datab1_add),     //   .datab
		.n         (n_add),         //   .n
		.reset     (reset),     //   .reset
		.reset_req (reset_req), //   .reset_req
		.start     (start_add),     //   .start
		.done      (done_add1),      //   .done
		.result    (result_add1)     //   .result
	);
	
fpoint2_multi #(
		.arithmetic_present (1),
		.root_present       (1),
		.conversion_present (1)
	) nios_custom_instr_floating_point_2_multi_2 (
		.clk       (clk),       // s1.clk
		.clk_en    (clk_en),    //   .clk_en
		.dataa     (dataa2_add),     //   .dataa
		.datab     (datab2_add),     //   .datab
		.n         (n_add),         //   .n
		.reset     (reset),     //   .reset
		.reset_req (reset_req), //   .reset_req
		.start     (start_add),     //   .start
		.done      (done_add2),      //   .done
		.result    (result_add2)     //   .result
	);
	
fpoint2_multi #(
		.arithmetic_present (1),
		.root_present       (1),
		.conversion_present (1)
	) nios_custom_instr_floating_point_2_multi_3 (
		.clk       (clk),       // s1.clk
		.clk_en    (clk_en),    //   .clk_en
		.dataa     (dataa3_add),     //   .dataa
		.datab     (datab3_add),     //   .datab
		.n         (n_add),         //   .n
		.reset     (reset),     //   .reset
		.reset_req (reset_req), //   .reset_req
		.start     (start_add),     //   .start
		.done      (done_add3),      //   .done
		.result    (result_add3)     //   .result
	);
	
fpoint2_multi #(
		.arithmetic_present (1),
		.root_present       (1),
		.conversion_present (1)
	) nios_custom_instr_floating_point_2_multi_4 (
		.clk       (clk),       // s1.clk
		.clk_en    (clk_en),    //   .clk_en
		.dataa     (dataa4_add),     //   .dataa
		.datab     (datab4_add),     //   .datab
		.n         (n_add),         //   .n
		.reset     (reset),     //   .reset
		.reset_req (reset_req), //   .reset_req
		.start     (start_add),     //   .start
		.done      (done_add4),      //   .done
		.result    (result_add4)     //   .result
	);

rise_edge_trigger ret1(
	.clk(clk),
	.reset(reset),
	.level(done_re_level),
	.rise_edge(next_in_edge)
);


hid_ram ramh(
	.address(address_hidden),
	.clock(clk),
	.data(wdata_hidden),
	.wren(wren_hidden),
	.q(rdata_hidden)
);

output_ram ramo(
	.address(address_out),
	.clock(clk),
	.data(wdata_out),
	.wren(wren_out),
	.q(rdata_out)
);



fp_max max(
	.clk(clk),
	.areset(reset),
	.a(dataa_comp),
	.b(datab_comp),
	.q(q_comp)
);



logic [31:0] wh1,wh2,wh3,wh4,rh1,rh2,rh3,rh4;
logic [31:0] wo1,wo2,ro1,ro2;
assign {wh4,wh3,wh2,wh1} = wdata_hidden;
assign {rh4,rh3,rh2,rh1} = rdata_hidden;
assign {wo2, wo1} = wdata_out;
assign {ro2, ro1} = rdata_out;


obs o1(
	.wh1(wh1),
	.wh2(wh2),
	.wh3(wh3),
	.wh4(wh4),
	.rh1(rh1),
	.rh2(rh2),
	.rh3(rh3),
	.rh4(rh4),
	.wo1(wo1),
	.wo2(wo2),
	.ro1(ro1),
	.ro2(ro2),
);

endmodule
