

module img_fifo (clk, reset, full, empty, wn, rn, datain, dataout);
  output reg [7:0] dataout;
  output full, empty;
  input [7:0] datain;
  input clk, reset, wn, rn;
  
  reg [9:0] wptr, rptr; // pointers tracking the stack
  reg [7:0] memory [783:0]; // the stack is 8 bit wide and 784 locations in size
  
  assign full = ( (wptr == 783) & (rptr == 0) ? 1 : 0 );
  assign empty = (wptr == rptr) ? 1 : 0;
  
  
  always @(posedge clk)
  begin
    if (reset)
      begin
        memory[0] <= 0;
memory[1] <= 0;
memory[2] <= 0;
memory[3] <= 0;
memory[4] <= 0;
memory[5] <= 0;
memory[6] <= 0;
memory[7] <= 0;
memory[8] <= 0;
memory[9] <= 0;
memory[10] <= 0;
memory[11] <= 0;
memory[12] <= 0;
memory[13] <= 0;
memory[14] <= 0;
memory[15] <= 0;
memory[16] <= 0;
memory[17] <= 0;
memory[18] <= 0;
memory[19] <= 0;
memory[20] <= 0;
memory[21] <= 0;
memory[22] <= 0;
memory[23] <= 0;
memory[24] <= 0;
memory[25] <= 0;
memory[26] <= 0;
memory[27] <= 0;
memory[28] <= 0;
memory[29] <= 0;
memory[30] <= 0;
memory[31] <= 0;
memory[32] <= 0;
memory[33] <= 0;
memory[34] <= 0;
memory[35] <= 0;
memory[36] <= 0;
memory[37] <= 0;
memory[38] <= 0;
memory[39] <= 0;
memory[40] <= 0;
memory[41] <= 0;
memory[42] <= 0;
memory[43] <= 0;
memory[44] <= 0;
memory[45] <= 0;
memory[46] <= 0;
memory[47] <= 0;
memory[48] <= 0;
memory[49] <= 0;
memory[50] <= 0;
memory[51] <= 0;
memory[52] <= 0;
memory[53] <= 0;
memory[54] <= 0;
memory[55] <= 0;
memory[56] <= 0;
memory[57] <= 0;
memory[58] <= 0;
memory[59] <= 0;
memory[60] <= 0;
memory[61] <= 0;
memory[62] <= 0;
memory[63] <= 0;
memory[64] <= 0;
memory[65] <= 0;
memory[66] <= 0;
memory[67] <= 0;
memory[68] <= 0;
memory[69] <= 0;
memory[70] <= 0;
memory[71] <= 0;
memory[72] <= 0;
memory[73] <= 0;
memory[74] <= 0;
memory[75] <= 0;
memory[76] <= 0;
memory[77] <= 0;
memory[78] <= 0;
memory[79] <= 0;
memory[80] <= 0;
memory[81] <= 0;
memory[82] <= 0;
memory[83] <= 0;
memory[84] <= 0;
memory[85] <= 0;
memory[86] <= 0;
memory[87] <= 0;
memory[88] <= 0;
memory[89] <= 0;
memory[90] <= 0;
memory[91] <= 0;
memory[92] <= 0;
memory[93] <= 0;
memory[94] <= 0;
memory[95] <= 0;
memory[96] <= 0;
memory[97] <= 0;
memory[98] <= 0;
memory[99] <= 0;
memory[100] <= 0;
memory[101] <= 0;
memory[102] <= 0;
memory[103] <= 0;
memory[104] <= 0;
memory[105] <= 0;
memory[106] <= 0;
memory[107] <= 0;
memory[108] <= 0;
memory[109] <= 0;
memory[110] <= 0;
memory[111] <= 0;
memory[112] <= 0;
memory[113] <= 0;
memory[114] <= 0;
memory[115] <= 0;
memory[116] <= 0;
memory[117] <= 0;
memory[118] <= 0;
memory[119] <= 0;
memory[120] <= 0;
memory[121] <= 0;
memory[122] <= 0;
memory[123] <= 0;
memory[124] <= 0;
memory[125] <= 0;
memory[126] <= 0;
memory[127] <= 0;
memory[128] <= 0;
memory[129] <= 0;
memory[130] <= 0;
memory[131] <= 0;
memory[132] <= 0;
memory[133] <= 0;
memory[134] <= 0;
memory[135] <= 0;
memory[136] <= 0;
memory[137] <= 0;
memory[138] <= 0;
memory[139] <= 0;
memory[140] <= 0;
memory[141] <= 0;
memory[142] <= 0;
memory[143] <= 0;
memory[144] <= 0;
memory[145] <= 0;
memory[146] <= 0;
memory[147] <= 0;
memory[148] <= 0;
memory[149] <= 0;
memory[150] <= 0;
memory[151] <= 0;
memory[152] <= 0;
memory[153] <= 0;
memory[154] <= 0;
memory[155] <= 0;
memory[156] <= 0;
memory[157] <= 0;
memory[158] <= 0;
memory[159] <= 0;
memory[160] <= 0;
memory[161] <= 0;
memory[162] <= 0;
memory[163] <= 0;
memory[164] <= 0;
memory[165] <= 0;
memory[166] <= 0;
memory[167] <= 0;
memory[168] <= 0;
memory[169] <= 0;
memory[170] <= 0;
memory[171] <= 0;
memory[172] <= 0;
memory[173] <= 0;
memory[174] <= 0;
memory[175] <= 0;
memory[176] <= 0;
memory[177] <= 0;
memory[178] <= 0;
memory[179] <= 0;
memory[180] <= 0;
memory[181] <= 0;
memory[182] <= 0;
memory[183] <= 0;
memory[184] <= 0;
memory[185] <= 0;
memory[186] <= 0;
memory[187] <= 0;
memory[188] <= 0;
memory[189] <= 0;
memory[190] <= 0;
memory[191] <= 0;
memory[192] <= 0;
memory[193] <= 0;
memory[194] <= 0;
memory[195] <= 0;
memory[196] <= 0;
memory[197] <= 0;
memory[198] <= 0;
memory[199] <= 0;
memory[200] <= 0;
memory[201] <= 0;
memory[202] <= 0;
memory[203] <= 0;
memory[204] <= 0;
memory[205] <= 0;
memory[206] <= 0;
memory[207] <= 0;
memory[208] <= 0;
memory[209] <= 0;
memory[210] <= 0;
memory[211] <= 0;
memory[212] <= 0;
memory[213] <= 0;
memory[214] <= 0;
memory[215] <= 0;
memory[216] <= 0;
memory[217] <= 0;
memory[218] <= 0;
memory[219] <= 0;
memory[220] <= 0;
memory[221] <= 0;
memory[222] <= 0;
memory[223] <= 0;
memory[224] <= 0;
memory[225] <= 0;
memory[226] <= 0;
memory[227] <= 0;
memory[228] <= 0;
memory[229] <= 0;
memory[230] <= 0;
memory[231] <= 0;
memory[232] <= 0;
memory[233] <= 0;
memory[234] <= 0;
memory[235] <= 0;
memory[236] <= 0;
memory[237] <= 0;
memory[238] <= 0;
memory[239] <= 0;
memory[240] <= 0;
memory[241] <= 0;
memory[242] <= 0;
memory[243] <= 0;
memory[244] <= 0;
memory[245] <= 0;
memory[246] <= 0;
memory[247] <= 0;
memory[248] <= 0;
memory[249] <= 0;
memory[250] <= 0;
memory[251] <= 0;
memory[252] <= 0;
memory[253] <= 0;
memory[254] <= 0;
memory[255] <= 0;
memory[256] <= 0;
memory[257] <= 0;
memory[258] <= 0;
memory[259] <= 0;
memory[260] <= 0;
memory[261] <= 0;
memory[262] <= 0;
memory[263] <= 0;
memory[264] <= 0;
memory[265] <= 0;
memory[266] <= 0;
memory[267] <= 0;
memory[268] <= 0;
memory[269] <= 0;
memory[270] <= 0;
memory[271] <= 0;
memory[272] <= 0;
memory[273] <= 0;
memory[274] <= 0;
memory[275] <= 0;
memory[276] <= 0;
memory[277] <= 0;
memory[278] <= 0;
memory[279] <= 0;
memory[280] <= 0;
memory[281] <= 0;
memory[282] <= 0;
memory[283] <= 0;
memory[284] <= 0;
memory[285] <= 0;
memory[286] <= 0;
memory[287] <= 0;
memory[288] <= 0;
memory[289] <= 0;
memory[290] <= 0;
memory[291] <= 0;
memory[292] <= 0;
memory[293] <= 0;
memory[294] <= 0;
memory[295] <= 0;
memory[296] <= 0;
memory[297] <= 0;
memory[298] <= 0;
memory[299] <= 0;
memory[300] <= 0;
memory[301] <= 0;
memory[302] <= 0;
memory[303] <= 0;
memory[304] <= 0;
memory[305] <= 0;
memory[306] <= 0;
memory[307] <= 0;
memory[308] <= 0;
memory[309] <= 0;
memory[310] <= 0;
memory[311] <= 0;
memory[312] <= 0;
memory[313] <= 0;
memory[314] <= 0;
memory[315] <= 0;
memory[316] <= 0;
memory[317] <= 0;
memory[318] <= 0;
memory[319] <= 0;
memory[320] <= 0;
memory[321] <= 0;
memory[322] <= 0;
memory[323] <= 0;
memory[324] <= 0;
memory[325] <= 0;
memory[326] <= 0;
memory[327] <= 0;
memory[328] <= 0;
memory[329] <= 0;
memory[330] <= 0;
memory[331] <= 0;
memory[332] <= 0;
memory[333] <= 0;
memory[334] <= 0;
memory[335] <= 0;
memory[336] <= 0;
memory[337] <= 0;
memory[338] <= 0;
memory[339] <= 0;
memory[340] <= 0;
memory[341] <= 0;
memory[342] <= 0;
memory[343] <= 0;
memory[344] <= 0;
memory[345] <= 0;
memory[346] <= 0;
memory[347] <= 0;
memory[348] <= 0;
memory[349] <= 0;
memory[350] <= 0;
memory[351] <= 0;
memory[352] <= 0;
memory[353] <= 0;
memory[354] <= 0;
memory[355] <= 0;
memory[356] <= 0;
memory[357] <= 0;
memory[358] <= 0;
memory[359] <= 0;
memory[360] <= 0;
memory[361] <= 0;
memory[362] <= 0;
memory[363] <= 0;
memory[364] <= 0;
memory[365] <= 0;
memory[366] <= 0;
memory[367] <= 0;
memory[368] <= 0;
memory[369] <= 0;
memory[370] <= 0;
memory[371] <= 0;
memory[372] <= 0;
memory[373] <= 0;
memory[374] <= 0;
memory[375] <= 0;
memory[376] <= 0;
memory[377] <= 0;
memory[378] <= 0;
memory[379] <= 0;
memory[380] <= 0;
memory[381] <= 0;
memory[382] <= 0;
memory[383] <= 0;
memory[384] <= 0;
memory[385] <= 0;
memory[386] <= 0;
memory[387] <= 0;
memory[388] <= 0;
memory[389] <= 0;
memory[390] <= 0;
memory[391] <= 0;
memory[392] <= 0;
memory[393] <= 0;
memory[394] <= 0;
memory[395] <= 0;
memory[396] <= 0;
memory[397] <= 0;
memory[398] <= 0;
memory[399] <= 0;
memory[400] <= 0;
memory[401] <= 0;
memory[402] <= 0;
memory[403] <= 0;
memory[404] <= 0;
memory[405] <= 0;
memory[406] <= 0;
memory[407] <= 0;
memory[408] <= 0;
memory[409] <= 0;
memory[410] <= 0;
memory[411] <= 0;
memory[412] <= 0;
memory[413] <= 0;
memory[414] <= 0;
memory[415] <= 0;
memory[416] <= 0;
memory[417] <= 0;
memory[418] <= 0;
memory[419] <= 0;
memory[420] <= 0;
memory[421] <= 0;
memory[422] <= 0;
memory[423] <= 0;
memory[424] <= 0;
memory[425] <= 0;
memory[426] <= 0;
memory[427] <= 0;
memory[428] <= 0;
memory[429] <= 0;
memory[430] <= 0;
memory[431] <= 0;
memory[432] <= 0;
memory[433] <= 0;
memory[434] <= 0;
memory[435] <= 0;
memory[436] <= 0;
memory[437] <= 0;
memory[438] <= 0;
memory[439] <= 0;
memory[440] <= 0;
memory[441] <= 0;
memory[442] <= 0;
memory[443] <= 0;
memory[444] <= 0;
memory[445] <= 0;
memory[446] <= 0;
memory[447] <= 0;
memory[448] <= 0;
memory[449] <= 0;
memory[450] <= 0;
memory[451] <= 0;
memory[452] <= 0;
memory[453] <= 0;
memory[454] <= 0;
memory[455] <= 0;
memory[456] <= 0;
memory[457] <= 0;
memory[458] <= 0;
memory[459] <= 0;
memory[460] <= 0;
memory[461] <= 0;
memory[462] <= 0;
memory[463] <= 0;
memory[464] <= 0;
memory[465] <= 0;
memory[466] <= 0;
memory[467] <= 0;
memory[468] <= 0;
memory[469] <= 0;
memory[470] <= 0;
memory[471] <= 0;
memory[472] <= 0;
memory[473] <= 0;
memory[474] <= 0;
memory[475] <= 0;
memory[476] <= 0;
memory[477] <= 0;
memory[478] <= 0;
memory[479] <= 0;
memory[480] <= 0;
memory[481] <= 0;
memory[482] <= 0;
memory[483] <= 0;
memory[484] <= 0;
memory[485] <= 0;
memory[486] <= 0;
memory[487] <= 0;
memory[488] <= 0;
memory[489] <= 0;
memory[490] <= 0;
memory[491] <= 0;
memory[492] <= 0;
memory[493] <= 0;
memory[494] <= 0;
memory[495] <= 0;
memory[496] <= 0;
memory[497] <= 0;
memory[498] <= 0;
memory[499] <= 0;
memory[500] <= 0;
memory[501] <= 0;
memory[502] <= 0;
memory[503] <= 0;
memory[504] <= 0;
memory[505] <= 0;
memory[506] <= 0;
memory[507] <= 0;
memory[508] <= 0;
memory[509] <= 0;
memory[510] <= 0;
memory[511] <= 0;
memory[512] <= 0;
memory[513] <= 0;
memory[514] <= 0;
memory[515] <= 0;
memory[516] <= 0;
memory[517] <= 0;
memory[518] <= 0;
memory[519] <= 0;
memory[520] <= 0;
memory[521] <= 0;
memory[522] <= 0;
memory[523] <= 0;
memory[524] <= 0;
memory[525] <= 0;
memory[526] <= 0;
memory[527] <= 0;
memory[528] <= 0;
memory[529] <= 0;
memory[530] <= 0;
memory[531] <= 0;
memory[532] <= 0;
memory[533] <= 0;
memory[534] <= 0;
memory[535] <= 0;
memory[536] <= 0;
memory[537] <= 0;
memory[538] <= 0;
memory[539] <= 0;
memory[540] <= 0;
memory[541] <= 0;
memory[542] <= 0;
memory[543] <= 0;
memory[544] <= 0;
memory[545] <= 0;
memory[546] <= 0;
memory[547] <= 0;
memory[548] <= 0;
memory[549] <= 0;
memory[550] <= 0;
memory[551] <= 0;
memory[552] <= 0;
memory[553] <= 0;
memory[554] <= 0;
memory[555] <= 0;
memory[556] <= 0;
memory[557] <= 0;
memory[558] <= 0;
memory[559] <= 0;
memory[560] <= 0;
memory[561] <= 0;
memory[562] <= 0;
memory[563] <= 0;
memory[564] <= 0;
memory[565] <= 0;
memory[566] <= 0;
memory[567] <= 0;
memory[568] <= 0;
memory[569] <= 0;
memory[570] <= 0;
memory[571] <= 0;
memory[572] <= 0;
memory[573] <= 0;
memory[574] <= 0;
memory[575] <= 0;
memory[576] <= 0;
memory[577] <= 0;
memory[578] <= 0;
memory[579] <= 0;
memory[580] <= 0;
memory[581] <= 0;
memory[582] <= 0;
memory[583] <= 0;
memory[584] <= 0;
memory[585] <= 0;
memory[586] <= 0;
memory[587] <= 0;
memory[588] <= 0;
memory[589] <= 0;
memory[590] <= 0;
memory[591] <= 0;
memory[592] <= 0;
memory[593] <= 0;
memory[594] <= 0;
memory[595] <= 0;
memory[596] <= 0;
memory[597] <= 0;
memory[598] <= 0;
memory[599] <= 0;
memory[600] <= 0;
memory[601] <= 0;
memory[602] <= 0;
memory[603] <= 0;
memory[604] <= 0;
memory[605] <= 0;
memory[606] <= 0;
memory[607] <= 0;
memory[608] <= 0;
memory[609] <= 0;
memory[610] <= 0;
memory[611] <= 0;
memory[612] <= 0;
memory[613] <= 0;
memory[614] <= 0;
memory[615] <= 0;
memory[616] <= 0;
memory[617] <= 0;
memory[618] <= 0;
memory[619] <= 0;
memory[620] <= 0;
memory[621] <= 0;
memory[622] <= 0;
memory[623] <= 0;
memory[624] <= 0;
memory[625] <= 0;
memory[626] <= 0;
memory[627] <= 0;
memory[628] <= 0;
memory[629] <= 0;
memory[630] <= 0;
memory[631] <= 0;
memory[632] <= 0;
memory[633] <= 0;
memory[634] <= 0;
memory[635] <= 0;
memory[636] <= 0;
memory[637] <= 0;
memory[638] <= 0;
memory[639] <= 0;
memory[640] <= 0;
memory[641] <= 0;
memory[642] <= 0;
memory[643] <= 0;
memory[644] <= 0;
memory[645] <= 0;
memory[646] <= 0;
memory[647] <= 0;
memory[648] <= 0;
memory[649] <= 0;
memory[650] <= 0;
memory[651] <= 0;
memory[652] <= 0;
memory[653] <= 0;
memory[654] <= 0;
memory[655] <= 0;
memory[656] <= 0;
memory[657] <= 0;
memory[658] <= 0;
memory[659] <= 0;
memory[660] <= 0;
memory[661] <= 0;
memory[662] <= 0;
memory[663] <= 0;
memory[664] <= 0;
memory[665] <= 0;
memory[666] <= 0;
memory[667] <= 0;
memory[668] <= 0;
memory[669] <= 0;
memory[670] <= 0;
memory[671] <= 0;
memory[672] <= 0;
memory[673] <= 0;
memory[674] <= 0;
memory[675] <= 0;
memory[676] <= 0;
memory[677] <= 0;
memory[678] <= 0;
memory[679] <= 0;
memory[680] <= 0;
memory[681] <= 0;
memory[682] <= 0;
memory[683] <= 0;
memory[684] <= 0;
memory[685] <= 0;
memory[686] <= 0;
memory[687] <= 0;
memory[688] <= 0;
memory[689] <= 0;
memory[690] <= 0;
memory[691] <= 0;
memory[692] <= 0;
memory[693] <= 0;
memory[694] <= 0;
memory[695] <= 0;
memory[696] <= 0;
memory[697] <= 0;
memory[698] <= 0;
memory[699] <= 0;
memory[700] <= 0;
memory[701] <= 0;
memory[702] <= 0;
memory[703] <= 0;
memory[704] <= 0;
memory[705] <= 0;
memory[706] <= 0;
memory[707] <= 0;
memory[708] <= 0;
memory[709] <= 0;
memory[710] <= 0;
memory[711] <= 0;
memory[712] <= 0;
memory[713] <= 0;
memory[714] <= 0;
memory[715] <= 0;
memory[716] <= 0;
memory[717] <= 0;
memory[718] <= 0;
memory[719] <= 0;
memory[720] <= 0;
memory[721] <= 0;
memory[722] <= 0;
memory[723] <= 0;
memory[724] <= 0;
memory[725] <= 0;
memory[726] <= 0;
memory[727] <= 0;
memory[728] <= 0;
memory[729] <= 0;
memory[730] <= 0;
memory[731] <= 0;
memory[732] <= 0;
memory[733] <= 0;
memory[734] <= 0;
memory[735] <= 0;
memory[736] <= 0;
memory[737] <= 0;
memory[738] <= 0;
memory[739] <= 0;
memory[740] <= 0;
memory[741] <= 0;
memory[742] <= 0;
memory[743] <= 0;
memory[744] <= 0;
memory[745] <= 0;
memory[746] <= 0;
memory[747] <= 0;
memory[748] <= 0;
memory[749] <= 0;
memory[750] <= 0;
memory[751] <= 0;
memory[752] <= 0;
memory[753] <= 0;
memory[754] <= 0;
memory[755] <= 0;
memory[756] <= 0;
memory[757] <= 0;
memory[758] <= 0;
memory[759] <= 0;
memory[760] <= 0;
memory[761] <= 0;
memory[762] <= 0;
memory[763] <= 0;
memory[764] <= 0;
memory[765] <= 0;
memory[766] <= 0;
memory[767] <= 0;
memory[768] <= 0;
memory[769] <= 0;
memory[770] <= 0;
memory[771] <= 0;
memory[772] <= 0;
memory[773] <= 0;
memory[774] <= 0;
memory[775] <= 0;
memory[776] <= 0;
memory[777] <= 0;
memory[778] <= 0;
memory[779] <= 0;
memory[780] <= 0;
memory[781] <= 0;
memory[782] <= 0;
memory[783] <= 0;

        dataout <= 0; wptr <= 0; rptr <= 0;
      end
    else if (wn & !full)
      begin
        memory[wptr] <= datain;
        wptr <= wptr + 1;
      end
    else if (rn & !empty)
      begin
        dataout <= memory[rptr];
        rptr <= rptr + 1;
      end
  end
endmodule